// Top Module 
module top(input wire clk12M,  // 12 MHz Clock pin (Lattice Board)
           input wire taster_reset, // Restart whole system and do sine stuff again
           output wire BLU);	  // Blue LED pin for onBoard LED (Lattice Board) 
  
  

  // Clocks
  wire sine_read_clk;  // Clock for generating 1MHz Sinewave
  wire clk_pwm; // need to be clk_read/resolution --> in our case: 1M/2^10 = 976.56 Hz
  wire clk24M;
  
  // Controll Signals
  wire write_finished;
  wire LED_PWM;
  wire valid;

  // Enable Signals 
  wire write_enable;
  wire read_enable;
  reg  enable_sin_gen_read;
  reg  enable_sin_write;

  // Reset Signals --> bring modules in defined states
  reg reset_RAM;
  reg reset_sin_gen;
  reg reset_write_sine;
  reg reset_pwm;
  
  // Data 
  wire [9:0] sine_val;
  wire [9:0] pwm_sin_val;
  wire [7:0] address_write;
  wire [7:0] address_read;
  wire [9:0] o_sin_value;
  wire LED_PWM;
  reg out_pwm;	
  
  
  PLL_24M PLL(.ref_clk_i(clk12M), 
			  .rst_n_i(reset_write_sine), 
			  .outcore_o(clk24M), 
			  .outglobal_o());
			  
  sine_gen SINGEN(.clk(sine_read_clk),
                  .enable(enable_sin_gen_read),
                  .address_read(address_read),
                  .data_sin_val(o_sin_value),
                  .pwm_sin_val(pwm_sin_val),
                  .reset(reset_sin_gen),
                  .data_valid(valid),
                  .read_enable(read_enable));
  

  write_sine SINWR(.clk(clk24M), 
                      .enable(enable_sin_write),
                  	  .reset(reset_write_sine),
                      .address_write(address_write),
                      .data_write(sine_val),
                      .write_finished(write_finished),
                      .write_enable(write_enable));
  
  pwm PWM(.clk(clk24M), .in_val(pwm_sin_val), .out_pwm(BLU), .enable(enable_sin_gen_read), .reset(reset_pwm), .valid(valid));
    
	
  RAM_LUT RAM(.wr_clk_i(clk24M), 
        .rd_clk_i(sine_read_clk), 
        .rst_i(reset_RAM), 
        .wr_clk_en_i(write_enable), 
        .rd_en_i(read_enable), 
        .rd_clk_en_i(read_enable), 
        .wr_en_i(write_enable), 
        .wr_data_i(sine_val), 
        .wr_addr_i(address_write), 
        .rd_addr_i(address_read), 
        .rd_data_o(o_sin_value));
		
  clock_devider  #(.WIDTH(12)) DIV(.reset(reset_pwm), .clk_in(clk24M), .clk_out(sine_read_clk)); // Generate 1/2^WIDTH of clk_in
  
  /* Dynamic behaviour:
  1. Step: Call Python Script to generate Sine Values
  2. Step: Reset Ram and enable write_sin module with "enable_sin_write"
  3. Step: Enable Sin_gen with enable_sin_gen_read
  	--> PWM Signal generated automatically by PWM Module 
  */
  
  initial begin
    // Reset RAM, sin_gen, sin_write, pwm  -> Reset whole System
    reset_RAM <= 1'b0;
  	reset_sin_gen <= 1'b0;
  	reset_write_sine <= 1'b0;
  	reset_pwm <= 1'b0;
    if(!reset_RAM) begin
      reset_RAM <= 1'b1;
      reset_sin_gen <= 1'b1;
      reset_write_sine <= 1'b1;
      reset_pwm <= 1'b1;
    end
    if(reset_RAM) begin
      reset_RAM <= 1'b0;
      reset_sin_gen <= 1'b0;
      reset_write_sine <= 1'b0;
      reset_pwm <= 1'b0;
    end
    
     enable_sin_gen_read = 1'b0;
 	 enable_sin_write = 1'b0;    
    
    // Fill RAM with values generated by Python Script
     enable_sin_write = 1'b1;
	 @(posedge write_finished)
      begin 
         enable_sin_write = 1'b0; // RAM filled
         enable_sin_gen_read = 1'b1; // Read RAM
      end
  end
  
  
  
  // uncomment and configure taster to add some additional functionallity
  // Restart Sine Generator at 
/*  always@(posedge taster_reset)begin

     enable_sin_gen_read = 1'b0; 
	 reset_sin_gen = 1'b1;
	 reset_pwm = 1'b1;
	 	
	if(reset_pwm) begin
		reset_sin_gen = 1'b0;  
		reset_pwm = 1'b0;
		enable_sin_write = 1'b1;    
	end
	
  end*/
  
  
endmodule
  