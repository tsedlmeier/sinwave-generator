// Moduel to write generated Sine values to RAM

module write_sine (clk, 
                  enable,				 
                  address_write,
                  data_write,
                  write_enable,
                  reset,
                  write_finished);
                  
input 			  clk;
input			  enable; 				 // enables whole module
input  			  reset;  
output  reg [7:0] address_write;
output  reg [9:0] data_write;
output  reg 	  write_enable;
output  reg		  write_finished;
integer i;
reg [9:0]  sine_vals [0:255];			// Array including Values of LUT

initial begin
  write_finished <= 1'b0;
  address_write <= 8'h00;
  data_write <= 10'b0000000000;
  write_enable <= 1'b0;
  i = 0;
  
  // Fill intern Array with write values : 
  // Path needs to be absolute 
  $readmemh("C:\\lscc\\radiant\\2.2\\projects\\sinewave_generator\\source\\impl_1\\ram_sine_vals.mem", sine_vals);
 end

  
  
 // Fill RAM with Sine Values
 // Values generated by python script
  always @(posedge clk ) begin  
	 if(reset) begin // Synchronous Reset
		address_write = 8'h00;
		data_write = 10'b0000000000;
		write_enable = 1'b0;   
		write_finished = 1'b0;
	end
    else if(enable) begin      	
        write_enable = 1'b1; 						// enables RAM write
        data_write = sine_vals[i];					// Write Value to RAM 
        address_write = address_write + 1'b1;       // Next address
    end
    
	if(address_write == 8'hFF) begin
      write_finished = 1'b1;						// Signals other Moduls that writing is finished now
      write_enable = 1'b0;
    end
    i = i +1;
  end
  

  
endmodule