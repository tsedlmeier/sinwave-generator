// Test Behaviour of submodules
`timescale 10ns/10ps
module test;
  
  wire sine_read_clk;
  reg clk;
  reg enable_sin_gen_read;
  reg enable_sin_write;
  wire write_finished;
  wire write_enable;
  wire read_enable;
  wire LED_PWM;
  wire valid;

  // Async Reset --> bring modules in defined states
  reg reset_RAM;
  reg reset_sin_gen;
  reg reset_write_sine;
  reg reset_pwm;
  
  wire [9:0] sine_val;
  wire [9:0] pwm_sin_val;
  wire [7:0] address_write;
  wire [7:0] address_read;
  wire [9:0] o_sin_value;

  sine_gen SINGEN(.clk(sine_read_clk),
                  .enable(enable_sin_gen_read),
                  .address_read(address_read),
                  .data_sin_val(o_sin_value),
                  .pwm_sin_val(pwm_sin_val),
                  .reset(reset_sin_gen),
                  .data_valid(valid),
                  .read_enable(read_enable));
  

  write_sine SINWR(.clk(clk), 
                      .enable(enable_sin_write),
                  	  .reset(reset_write_sine),
                      .address_write(address_write),
                      .data_write(sine_val),
                      .write_finished(write_finished),
                      .write_enable(write_enable));
  
  pwm PWM(.clk(clk), .in_val(pwm_sin_val), .out_pwm(LED_PWM), .enable(enable_sin_gen_read), .reset(reset_pwm), .valid(valid));
  

  RAM_LUT RAM(.wr_clk_i(clk), 
        .rd_clk_i(sine_read_clk), 
        .rst_i(reset_RAM), 
        .wr_clk_en_i(write_enable), 
        .rd_en_i(read_enable), 
        .rd_clk_en_i(read_enable), 
        .wr_en_i(write_enable), 
        .wr_data_i(sine_val), 
        .wr_addr_i(address_write), 
        .rd_addr_i(address_read), 
        .rd_data_o(o_sin_value));
		
  clock_devider #(.WIDTH(10)) DIV(.reset(reset_pwm), .clk_in(clk), .clk_out(sine_read_clk));
  
  initial begin

    clk = 1'b0;
	//clk24M = 1'b0;
	//sine_read_clk = 1'b0;
    
    // Reset RAM, sin_gen, sin_write, pwm  -> Reset whole System
    reset_RAM <= 1'b0;
  	reset_sin_gen <= 1'b0;
  	reset_write_sine <= 1'b0;
  	reset_pwm <= 1'b0;
    if(!reset_RAM) begin
      reset_RAM <= 1'b1;
      reset_sin_gen <= 1'b1;
      reset_write_sine <= 1'b1;
      reset_pwm <= 1'b1;
    end
    if(reset_RAM) begin
      reset_RAM <= 1'b0;
      reset_sin_gen <= 1'b0;
      reset_write_sine <= 1'b0;
      reset_pwm <= 1'b0;
    end
    
     enable_sin_gen_read = 1'b0;
 	 enable_sin_write = 1'b0;    
    
    // Fill RAM with values generated by Python Script
     enable_sin_write = 1'b1;
	 @(posedge write_finished)
      begin 
         enable_sin_write = 1'b0; // RAM filled
         enable_sin_gen_read = 1'b1; // Read RAM
      end
 end
    
    

  // Generate Clocks
  always #8.3 clk = ~clk; // 12 MHz Clock from board
  //always #8.3 clk = ~clk; // 12 MHz Clock from board
  //always #8.3 clk = ~clk; // 12 MHz Clock from board
  
endmodule